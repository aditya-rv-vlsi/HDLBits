module top_module ( input [1:0] A, input [1:0] B, output z ); 
    z = (A==B)?1:0;
endmodule
